`timescale 1ns / 1ps

module InstructionMem(
    input [31:0] inport1,
    input readIM,
    output reg [31:0] R1
);
    reg [31:0] R[255:0];
    
    initial begin
    //    R[0] = 32'b11000000000000000000000000000010;//BR 2
    //    R[0] = 32'b01000110000000000000000001100001;//BPL R6,3
    //    R[1] = 32'b00000001000000010100000000000000;
    //    R[2] = 32'b00100011001010000000000000100001;
    //    R[3] = 32'b00100011000010000000000000000000;
    //     R[4] = 32'b00100011000100000000000000100000;
    //    R[5] = 32'b00000001000100010000000000001000;//ADD R4,R1.R2
    //    R[6] = 32'b01000000000111111111111100100011;

        // gcd
        R[0]=32'b00000001000100010000000000000010;
        R[1]=32'b01000100000000000000000010100011;
        R[2]=32'b01000100000000000000000001000001;
        R[3]=32'b00000001000100000100000000000010;
        R[4]=32'b11000011111111111111111111111011;
        R[5]=32'b00000010000010001000000000000010;
        R[6]=32'b11000011111111111111111111111001;
        R[7]=32'b00000001000000001100000000000000;
        R[8]=32'b11000011111111111111111111111111;

        //booth
        // R[0] = 32'b00000000000000010100000000000000;
        // R[1] = 32'b00000000000000011000000000000000;
        // R[2] = 32'b00000000000000011100000000000000;
        // R[3] = 32'b00000111000000000000000111100001;
        // R[4] = 32'b01000111000000000000001011000011;
        // R[5] = 32'b00000010000000100000000000000000;
        // R[6] = 32'b00001000000000000000000000100101;
        // R[7] = 32'b01001000000000000000000001000011;
        // R[8] = 32'b01000110000000000000000010000011;
        // R[9] = 32'b11000000000000000000000000000100;
        // R[10] = 32'b01000110000000000000000001100011;
        // R[11] = 32'b00000101000010010100000000000000;
        // R[12] = 32'b11000000000000000000000000000001;
        // R[13] = 32'b00000101000010010100000000000010;
        // R[14] = 32'b00000000000000011000000000000000;
        // R[15] = 32'b01001000000000000000000000100011;
        // R[16] = 32'b00000110000000000000000000100001;
        // R[17] = 32'b00000010000000000000000000101110;
        // R[18] = 32'b00000101000000100000000000000000;
        // R[19] = 32'b00001000000000000000000000100101;
        // R[20] = 32'b01001000000000000000000001000011;
        // R[21] = 32'b00000010000010000000000000000111;
        // R[22] = 32'b11000000000000000000000000000001;
        // R[23] = 32'b00000010000001111111111111100101;
        // R[24] = 32'b00000101000000000000000000101110;
        // R[25] = 32'b00000111000000000000000000100011;
        // R[26] = 32'b11000011111111111111111111101001;
        // R[27] = 32'b00000101000000001100000000000000;
        // R[28] = 32'b00000010000000010000000000000000;
        // R[29] = 32'b11000011111111111111111111111111;
    end
    
    always @(*) begin
        if(readIM == 1'b1)
        R1=R[inport1];
    end
endmodule

